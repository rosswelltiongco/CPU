`timescale 1ns / 1ps
/********************************************************************************
 *
 * Author:   Rosswell Tiongco & Jesus Luciano
 * Email:    rosswelltiongco@gmail.com & jlucian995@gmail.com
 * Filename: top_level_lab5.v
 * Date:     
 * Version:  1.0
 *
 * Description: 
 *
 *
 *******************************************************************************/
module top_level_lab5();


endmodule
