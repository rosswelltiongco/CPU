`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:31:55 10/11/2017 
// Design Name: 
// Module Name:    pixel_controller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module pixel_controller(
    input clk,
    input reset,
    output a7,
    output a6,
    output a5,
    output a4,
    output a3,
    output a2,
    output a1,
    output a0,
    output [2:0] seg_sel
    );


endmodule
