`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:30:47 10/11/2017 
// Design Name: 
// Module Name:    ad_mux 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ad_mux(
    input [3:0] d7,
    input [3:0] d6,
    input [3:0] d5,
    input [3:0] d4,
    input [3:0] d3,
    input [3:0] d2,
    input [3:0] d1,
    input [3:0] d0,
    input [2:0] sel,
    output [3:0] Y
    );


endmodule
